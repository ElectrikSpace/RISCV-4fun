ROM_block_inst : ROM_block PORT MAP (
		address_a	 => address_a_sig,
		address_b	 => address_b_sig,
		clock_a	 => clock_a_sig,
		clock_b	 => clock_b_sig,
		enable_a	 => enable_a_sig,
		enable_b	 => enable_b_sig,
		q_a	 => q_a_sig,
		q_b	 => q_b_sig
	);
